module Final_Project(clk, rst, button, VGA_CLK, VGA_VS, VGA_HS, VGA_BLANK_N, VGA_SYNC_N, VGA_R, VGA_G, VGA_B, light1, light2, seg7_neg_sign, seg7_digmsb, seg7_digmid, seg7_diglsb);
	input clk;
	input rst;
	input [1:0] button;

	// Outputs used by the VGA module.
	output VGA_CLK;
	output VGA_HS;
	output VGA_VS;
	output VGA_BLANK_N;
	output VGA_SYNC_N;
	output [9:0] VGA_R;
	output [9:0] VGA_G;
	output [9:0] VGA_B;
	
	// Used for quick debugging.
	output reg light1;
	output reg light2;
	
	output [6:0]seg7_neg_sign;
	output [6:0]seg7_digmsb;
	output [6:0]seg7_digmid;
	output [6:0]seg7_diglsb;

	// Instantiate the VGA module (received from previous students of 287).
	vga_adapter VGA(
	  .resetn(1'b1),
	  .clock(clk),
	  .colour(colour),
	  .x(x),
	  .y(y),
	  .plot(1'b1),
	  .VGA_R(VGA_R),
	  .VGA_G(VGA_G),
	  .VGA_B(VGA_B),
	  .VGA_HS(VGA_HS),
	  .VGA_VS(VGA_VS),
	  .VGA_BLANK(VGA_BLANK_N),
	  .VGA_SYNC(VGA_SYNC_N),
	  .VGA_CLK(VGA_CLK));
	defparam VGA.RESOLUTION = "160x120";
	defparam VGA.MONOCHROME = "FALSE";
	defparam VGA.BITS_PER_COLOUR_CHANNEL = 2;
	defparam VGA.BACKGROUND_IMAGE = "";
	
	clock frameKeeper(.clock(clk), .clk(frame));
	two_decimal_vals_w_neg splitter(player_balance, seg7_neg_sign, seg7_diglsb, seg7_digmid, seg7_digmsb);
	
	
	reg [9:0]player_balance;
	reg [7:0]S;
	reg [7:0]NS;
	reg [17:0]draw;
	reg done;
	reg spinReady;
	
	reg [7:0]x;
	reg [7:0]y;
	reg [5:0]colour;
	
	wire frame;
	wire [2:0]rand1;
	wire [2:0]rand2;
	wire [2:0]rand3;
	

	parameter backgroundImageBits = 4096'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000001000000000000000000000000000000000000000001000000000000000000000000000000000000000000001100000000000000000000000000000000000000010000000000000000000000000000000000000000010000000000000000000000000000000000000000000011000000000000000000000000000000000000000100000000000000000000000000000000000000000100000000000000000000000000000000000000000000110000000000000000000000000000000000000001000000000000000000000000000000000000000001000000000000000000000000000000000000000000001100000000000000000000000000000000000000010000000000000000000000000000000000000000010000000000000000000000000000000000000000000011000000000000000000000000000000000000000100000000000000000000000000000000000000000100000000000000000000000000000000000000000000110000000000000000000000000000000000000001000000000000000000000000000000000000000001000000000000000000000000000000000000000000001100000000000000000000000000000000000000010000000000000000000000000000000000000000010000000000000000000000000000000000000000000011000000000000000000000000000000000000000100000000000000000000000000000000000000000100000000000000000000000000000000000000000000110000000000000000000000000000000000000001000000000000000000000000000000000000000001000000000000000000000000000000000000000000001100000000000000000000000000000000000000010000000000000000000000000000000000000000010000000000000000000000000000000000000000000011000000000000000000000000000000000000000100000000000000000000000000000000000000000100000000000000000000000000000000000000000000110000000000000000000000000000000000000001000000000000000000000000000000000000000001000000000000000000000000000000000000000000001100000000000000000000000000000000000000010000000000000000000000000000000000000000010000000000000000000000000000000000000000000011000000000000000000000000000000000000000100000000000000000000000000000000000000000100000000000000000000000000000000000000000000110000000000000000000000000000000000000001000000000000000000000000000000000000000001000000000000000000000000000000000000000000001100000000000000000000000000000000000000010000000000000000000000000000000000000000010000000000000000000000000000000000000000000011000000000000000000000000000000000000000100000000000000000000000000000000000000000100000000000000000000000000000000000000000000110000000000000000000000000000000000000001000000000000000000000000000000000000000001000000000000000000000000000000000000000000001100000000000000000000000000000000000000010000000000000000000000000000000000000000010000000000000000000000000000000000000000000011000000000000000000000000000000000000000100000000000000000000000000000000000000000100000000000000000000000000000000000000000000110000000000000000000000000000000000000001000000000000000000000000000000000000000001000000000000000000000000000000000000000000001100000000000000000000000000000000000000010000000000000000000000000000000000000000010000000000000000000000000000000000000000000011000000000000000000000000000000000000000100000000000000000000000000000000000000000100000000000000000000000000000000000000000000110000000000000000000000000000000000000001000000000000000000000000000000000000000001000000000000000000000000000000000000000000001100000000000000000000000000000000000000010000000000000000000000000000000000000000010000000000000000000000000000000000000000000011000000000000000000000000000000000000000100000000000000000000000000000000000000000100000000000000000000000000000000000000000000110000000000000000000000000000000000000001000000000000000000000000000000000000000001000000000000000000000000000000000000000000001100000000000000000000000000000000000000010000000000000000000000000000000000000000010000000000000000000000000000000000000000000011000000000000000000000000000000000000000100000000000000000000000000000000000000000100000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
				 backgroundImageWidth = 63'd127,
				 backgroundImageHeight = 7'd32,
				 backgroundImageStart = 12'd4095;
				 
	parameter winImageBits = 4096'b0000000000000000111100000000000000011110000000000000000111100000011110000000000111100000000000000001110000000000000000000000000000000000000000001111000000000000000111110000000000000011111000000111100000000011111110000000000000011110000000000000000000000000000000000000000011111000000000000011111100000000000000111110000001111000000000111111110000000000000111100000000000000000000000000000000000000000111110000000000000111111000000000000001111000000011110000000001111111100000000000001111000000000000000000000000000000000000000000111100000000000001111111000000000000011110000000111100000000011111111100000000000011110000000000000000000000000000000000000000001111100000000000011111110000000000001111100000001111000000000111111111000000000000111100000000000000000000000000000000000000000011111000000000001111111100000000000011111000000011110000000001111011111000000000001111000000000000000000000000000000000000000000111110000000000011111111000000000000111100000000111100000000011110011110000000000011110000000000000000000000000000000000000000000111100000000000111111111000000000001111000000001111000000000111100111110000000000111100000000000000000000000000000000000000000001111100000000001111011110000000000111110000000011110000000001111000111100000000001111000000000000000000000000000000000000000000011111000000000111100111100000000001111000000000111100000000011111001111100000000011110000000000000000000000000000000000000000000011110000000001111001111100000000011110000000001111000000000111110001111000000000111100000000000000000000000000000000000000000000111100000000011110011111000000000111100000000011110000000001111100011111000000001111000000000000000000000000000000000000000000001111100000000111100011110000000011111000000000111100000000011111000011111000000011110000000000000000000000000000000000000000000001111000000011110000111100000000111100000000001111000000000111110000111110000000111100000000000000000000000000000000000000000000011110000000111100001111100000001111000000000011110000000001111100000111110000001111000000000000000000000000000000000000000000000111100000001111000001111000000011110000000000111100000000011111000001111100000011110000000000000000000000000000000000000000000001111100000011100000011110000001111000000000001111000000000111110000001111100000111100000000000000000000000000000000000000000000001111000001111000000111100000011110000000000011110000000001111100000011111000001111000000000000000000000000000000000000000000000011110000011110000001111100000111100000000000111100000000011111000000011111000011110000000000000000000000000000000000000000000000111110000111100000001111000011110000000000001111000000000111110000000111110000111100000000000000000000000000000000000000000000000111100001110000000011110000111100000000000011110000000001111100000000111110001111000000000000000000000000000000000000000000000001111000111100000000111110001111000000000000111100000000011111000000000111100011110000000000000000000000000000000000000000000000011110001111000000000111100011110000000000001111000000000111110000000001111100111100000000000000000000000000000000000000000000000111110011110000000001111001111000000000000011110000000001111100000000001111001111000000000000000000000000000000000000000000000000111100111000000000011110011110000000000000111100000000011111000000000011111011110000000000000000000000000000000000000000000000001111011110000000000111110111100000000000001111000000000111110000000000011111111100000000000000000000000000000000000000000000000011110111100000000000111101110000000000000011110000000001111100000000000111111111000000000000000000000000000000000000000000000000011111111000000000001111111100000000000000111100000000011111000000000000111111110000000000000000000000000000000000000000000000000111111100000000000011111111000000000000001111000000000111110000000000001111111100000000000000000000000000000000000000000000000001111111000000000000011111110000000000000011110000000001111100000000000001111111000000000000000000000000000000000000000000000000011111110000000000000111111000000000000000111100000000011111000000000000011111110000000000000000000000000,
				 winImageWidth = 63'd127,
				 winImageHeight = 7'd32,
				 winImageStart = 12'd4095;
				 
	parameter loseImageBits = 4096'b0000000000000000111100000000000000000000000001111111111100000000000000000001111111110000000000001111111111111111000000000000000000000000000000001111000000000000000000000001111111111111110000000000000001111111111111000000000111111111111111111000000000000000000000000000000011110000000000000000000001111111111111111110000000000000111111111111111000000001111111111111111110000000000000000000000000000000111100000000000000000000111111111001111111111000000000011111110001111110000000011111111111111111000000000000000000000000000000001111000000000000000000011111100000000001111110000000001111110000000011100000000111100000000000000000000000000000000000000000000011110000000000000000001111110000000000001111110000000011111000000000000000000001111000000000000000000000000000000000000000000000111100000000000000000011111000000000000001111110000000111100000000000000000000011110000000000000000000000000000000000000000000001111000000000000000001111100000000000000001111100000001111000000000000000000000111100000000000000000000000000000000000000000000011110000000000000000011111000000000000000001111000000011110000000000000000000001111000000000000000000000000000000000000000000000111100000000000000001111100000000000000000011111000000111100000000000000000000011110000000000000000000000000000000000000000000001111000000000000000011111000000000000000000111110000001111100000000000000000000111100000000000000000000000000000000000000000000011110000000000000000111110000000000000000000111100000011111100000000000000000001111000000000000000000000000000000000000000000000111100000000000000001111000000000000000000001111000000011111100000000000000000011110000000000000000000000000000000000000000000001111000000000000000011110000000000000000000011110000000111111110000000000000000111100000000000000000000000000000000000000000000011110000000000000000111100000000000000000000111110000000111111111000000000000001111111111111111000000000000000000000000000000000111100000000000000001111000000000000000000001111100000000011111111100000000000011111111111111110000000000000000000000000000000001111000000000000000011110000000000000000000011111000000000011111111110000000000111111111111111100000000000000000000000000000000011110000000000000000111100000000000000000000111110000000000001111111110000000001111100000000000000000000000000000000000000000000111100000000000000001111000000000000000000001111000000000000000011111110000000011110000000000000000000000000000000000000000000001111000000000000000011110000000000000000000011110000000000000000011111110000000111100000000000000000000000000000000000000000000011110000000000000000111100000000000000000000111100000000000000000001111100000001111000000000000000000000000000000000000000000000111100000000000000001111100000000000000000011111000000000000000000001111100000011110000000000000000000000000000000000000000000001111000000000000000011111000000000000000000111110000000000000000000011111000000111100000000000000000000000000000000000000000000011110000000000000000111110000000000000000001111000000000000000000000111110000001111000000000000000000000000000000000000000000000111100000000000000000111110000000000000000111110000000000000000000001111100000011110000000000000000000000000000000000000000000001111000000000000000001111100000000000000001111100000000000000000000011111000000111100000000000000000000000000000000000000000000011110000000000000000011111100000000000000111110000000000000000000000111100000001111000000000000000000000000000000000000000000000111100000000000000000011111100000000000011111100000001100000000000011111000000011110000000000000000000000000000000000000000000001111000000000000000000011111110000000011111110000000011110000000001111100000000111100000000000000000000000000000000000000000000011111111111111110000000011111111111111111111000000000111111111111111111000000001111111111111111110000000000000000000000000000000111111111111111110000000011111111111111111100000000001111111111111111100000000011111111111111111100000000000000000000000000000001111111111111111000000000011111111111111100000000000000111111111111100000000000111111111111111111000000000000000,
				 loseImageWidth = 63'd127,
				 loseImageHeight = 7'd32,
				 loseImageStart = 12'd4095;
	
	parameter startImageBits = 512'b00000000000000000000000000000000001111111111111001111111111111000011111111111110011111111111110000111100000000000110000000001100001111000000000001100000000011000011110000000000011000000000110000111100000011100110000000001100001111000000111001100000000011000011110000000110011000000000110000111111111111100111111111111100001111111111111001111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	          startImageWidth = 5'd31,
				 startImageHeight = 5'd16,
				 startImageStart = 9'd511;
				 
	parameter sevenImageBits = 512'b00000000000000000000000000000000000001111111111111111111111000000000011111111111111111111110000000000111111111111111111111100000000000000000000000111111111000000000000000000000011111111100000000000000000000001111111110000000000000000000000111111111000000000000000000000011111111100000000000000000000001111111110000000000000000000000111111111000000000000000000000011111111100000000000000000000001111111110000000000000000000000111111111000000000000000000000011111111100000000000000000000000000000000000000000000000,
				 sevenImageWidth = 5'd31,
				 sevenImageHeight = 5'd16,
				 sevenImageStart = 9'd511;
				 
	parameter orangeImageBits = 512'b00000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000001111111111111100000000000000000111111111111111100000000000000011111111111111111100000000000001111111111111111111100000000000111111111111111111111100000000000111111111111111111110000000000000111111111111111111000000000000000111111111111111100000000000000000111111111111110000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
				 orangeImageWidth = 5'd31,
				 orangeImageHeight = 5'd16,
				 orangeImageStart = 9'd511;
				 
	parameter lemonImageBits = 512'b00000000000000000000000000000000000000000000011110000000000000000000000000011111111000000000000000000000001111111111000000000000000000000111111111111000000000000000000011111111111111000000000000000001111111111111111000000000000000011111111111111110000000000000000011111111111111000000000000000000011111111111100000000000000000000011111111110000000000000000000000011111111000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
				 lemonImageWidth = 5'd31,
				 lemonImageHeight = 5'd16,
				 lemonImageStart = 9'd511;
				 
	parameter coinImageBits = 512'b00000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000001000000100000100000000000000000100111111111100100000000000000010001100010000000100000000000001000011000100000000100000000000100000110001000000000100000000000100001100010000000010000000000000100011000100000001000000000000000100111111111100100000000000000000100000010000010000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
				 coinImageWidth = 5'd31,
				 coinImageHeight = 5'd16,
				 coinImageStart = 9'd511;
				 
	parameter dollarImageBits = 512'b00000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000000000000001111111111111111110000000000000010000000010000000000000000000000100000000100000000000000000000001000000001000000000000000000000010000000010000000000000000000000111111111111111111000000000000000000000001000000010000000000000000000000010000000100000000000000000000000100000001000000000000000000000001000000010000000000000011111111111111111100000000000000000000000100000000000000000000000000000001000000000000000,
				 dollarImageWidth = 5'd31,
				 dollarImageHeight = 5'd16,
				 dollarImageStart = 9'd511;
				 
	parameter boltImageBits = 512'b00000000000000000000000000000000000000001000000000000000111100000000000000000000000000111100000000001000000000000000111110000000000000000000000000011111100000000000000000000000001111110000000000000001000000111111010000000000000000000001111111110000001000000000000000111111111000000000000000000000011111100000010000000000000000001111100000000000000000000000000011111000000000000000000000000011111000000010000000100000000001111100000000000000000000000001111100000000000000000000000000000000000000000000000000000000,
				 boltImageWidth = 5'd31,
				 boltImageHeight = 5'd16,
				 boltImageStart = 9'd511;
				 
	parameter bombImageBits = 512'b00000000000000000000000000000000000000001110000000000000000000000000000001110000000000000000000000000000001110000000000000000000000000001111111111110000000000000000000111111111111110000000000000000011111111111111110000000000000001111111111111111110000000000000111111111111111111110000000000011111111111111111111110000000000011111111111111111111000000000000011111111111111111100000000000000011111111111111110000000000000000011111111111111000000000000000000011111111111100000000000000000000000000000000000000000000,
				 bombImageWidth = 5'd31,
				 bombImageHeight = 5'd16,
				 bombImageStart = 9'd511;
				 
	parameter clearImageBits = 512'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
				 clearImageWidth = 5'd31,
				 clearImageHeight = 5'd16,
				 clearImageStart = 9'd511;

				 
	reg [63:0]imageX;
	reg [63:0]imageY;
	reg [63:0]counter;
	reg [63:0]currentInitX;
	reg [2:0]currentLeftSlot;
	reg [2:0]currentMidSlot;
	reg [2:0]currentRightSlot;
	reg [1:0]currentCheckState;
	reg [63:0]debounceCounter;
	reg [4:0]loopCounter;
	
	parameter initXBG = 63'd15,
			    initYBG = 63'd15,
				 initXStartLeftSlot = 63'd19,
				 initYStartLeftSlot = 63'd22,
				 initXStartMidSlot = 63'd60,
				 initYStartMidSlot = 63'd22,
				 initXStartRightSlot = 63'd103,
				 initYStartRightSlot = 63'd22,
				 initXEnd = 63'd15,
				 initYEnd = 63'd55;
	
	parameter START = 8'd0,
				 START_DRAW_BG = 8'd1,
				 INIT_DRAW_BG = 8'd2,
				 COND_DRAW_BG = 8'd3,
				 DRAW_BG = 8'd4,
				 BITCOND_DRAW_BG = 8'd5,
				 INCX_DRAW_BG = 8'd6,
				 INCY_DRAW_BG = 8'd7,
				 DEC_COUNTER_DRAW_BG = 8'd8,
				 EXIT_DRAW_BG = 8'd9,
				 
				 
				 init_left_slot = 8'd10,
				 START_DRAW_START_LEFT = 8'd11,
				 INIT_DRAW_START_LEFT = 8'd12,
				 COND_DRAW_START_LEFT = 8'd13,
				 DRAW_START_LEFT = 8'd14,
				 BITCOND_DRAW_START_LEFT = 8'd15,
				 INCX_DRAW_START_LEFT = 8'd16,
				 INCY_DRAW_START_LEFT = 8'd17,
				 DEC_COUNTER_DRAW_START_LEFT = 8'd18,
				 EXIT_DRAW_START_LEFT = 8'd19,
				 
				 
				 init_mid_slot = 8'd20,
				 START_DRAW_START_MID = 8'd21,
				 INIT_DRAW_START_MID = 8'd22,
				 COND_DRAW_START_MID = 8'd23,
				 DRAW_START_MID = 8'd24,
				 BITCOND_DRAW_START_MID = 8'd25,
				 INCX_DRAW_START_MID = 8'd26,
				 INCY_DRAW_START_MID = 8'd27,
				 DEC_COUNTER_DRAW_START_MID = 8'd28,
				 EXIT_DRAW_START_MID = 8'd29,
				 
				 
				 init_right_slot = 8'd30,
				 START_DRAW_START_RIGHT = 8'd31,
				 INIT_DRAW_START_RIGHT = 8'd32,
				 COND_DRAW_START_RIGHT = 8'd33,
				 DRAW_START_RIGHT = 8'd34,
				 BITCOND_DRAW_START_RIGHT = 8'd35,
				 INCX_DRAW_START_RIGHT = 8'd36,
				 INCY_DRAW_START_RIGHT = 8'd37,
				 DEC_COUNTER_DRAW_START_RIGHT = 8'd38,
				 EXIT_DRAW_START_RIGHT = 8'd39,
				 
				 CLEAR_SLOTS = 8'd40,
				 
				 START_CLEAR_LEFT = 8'd41,
				 INIT_CLEAR_LEFT = 8'd42,
				 COND_CLEAR_LEFT = 8'd43,
				 CLEAR_LEFT = 8'd44,
				 BITCOND_CLEAR_LEFT = 8'd45,
				 INCX_CLEAR_LEFT = 8'd46,
				 INCY_CLEAR_LEFT = 8'd47,
				 DEC_COUNTER_CLEAR_LEFT = 8'd48,
				 EXIT_CLEAR_LEFT = 8'd49,
				 
				 START_CLEAR_MID = 8'd50,
				 INIT_CLEAR_MID = 8'd51,
				 COND_CLEAR_MID = 8'd52,
				 CLEAR_MID = 8'd53,
				 BITCOND_CLEAR_MID = 8'd54,
				 INCX_CLEAR_MID = 8'd55,
				 INCY_CLEAR_MID = 8'd56,
				 DEC_COUNTER_CLEAR_MID = 8'd57,
				 EXIT_CLEAR_MID = 8'd58,
				 
				 START_CLEAR_RIGHT = 8'd59,
				 INIT_CLEAR_RIGHT = 8'd60,
				 COND_CLEAR_RIGHT = 8'd61,
				 CLEAR_RIGHT = 8'd62,
				 BITCOND_CLEAR_RIGHT = 8'd63,
				 INCX_CLEAR_RIGHT = 8'd64,
				 INCY_CLEAR_RIGHT = 8'd65,
				 DEC_COUNTER_CLEAR_RIGHT = 8'd66,
				 EXIT_CLEAR_RIGHT = 8'd67,
				 
				 WAIT_FOR_INPUT = 8'd68,
				 CHECK_SLOT1 = 8'd69,
				 CHECK_SLOT2 = 8'd70,
				 CHECK_SLOT3 = 8'd71,
				 
				 START_DRAW_SEVEN = 8'd72,
				 INIT_DRAW_SEVEN = 8'd73,
				 COND_DRAW_SEVEN = 8'd74,
				 DRAW_SEVEN = 8'd75,
				 BITCOND_DRAW_SEVEN = 8'd76,
				 INCX_DRAW_SEVEN = 8'd77,
				 INCY_DRAW_SEVEN = 8'd78,
				 DEC_COUNTER_DRAW_SEVEN = 8'd79,
				 EXIT_DRAW_SEVEN = 8'd80,
				 
				 START_DRAW_ORANGE = 8'd81,
				 INIT_DRAW_ORANGE = 8'd82,
				 COND_DRAW_ORANGE = 8'd83,
				 DRAW_ORANGE = 8'd84,
				 BITCOND_DRAW_ORANGE = 8'd85,
				 INCX_DRAW_ORANGE = 8'd86,
				 INCY_DRAW_ORANGE = 8'd87,
				 DEC_COUNTER_DRAW_ORANGE = 8'd88,
				 EXIT_DRAW_ORANGE = 8'd89,
				 
				 START_DRAW_LEMON = 8'd90,
				 INIT_DRAW_LEMON = 8'd91,
				 COND_DRAW_LEMON = 8'd92,
				 DRAW_LEMON = 8'd93,
				 BITCOND_DRAW_LEMON = 8'd94,
				 INCX_DRAW_LEMON = 8'd95,
				 INCY_DRAW_LEMON = 8'd96,
				 DEC_COUNTER_DRAW_LEMON = 8'd97,
				 EXIT_DRAW_LEMON = 8'd98,
				 
				 START_DRAW_COIN = 8'd99,
				 INIT_DRAW_COIN = 8'd100,
				 COND_DRAW_COIN = 8'd101,
				 DRAW_COIN = 8'd102,
				 BITCOND_DRAW_COIN = 8'd103,
				 INCX_DRAW_COIN = 8'd104,
				 INCY_DRAW_COIN = 8'd105,
				 DEC_COUNTER_DRAW_COIN = 8'd106,
				 EXIT_DRAW_COIN = 8'd107,
				 
				 START_DRAW_DOLLAR = 8'd108,
				 INIT_DRAW_DOLLAR = 8'd109,
				 COND_DRAW_DOLLAR = 8'd110,
				 DRAW_DOLLAR = 8'd111,
				 BITCOND_DRAW_DOLLAR = 8'd112,
				 INCX_DRAW_DOLLAR = 8'd113,
				 INCY_DRAW_DOLLAR = 8'd114,
				 DEC_COUNTER_DRAW_DOLLAR = 8'd115,
				 EXIT_DRAW_DOLLAR = 8'd116,
				 
				 START_DRAW_BOLT = 8'd117,
				 INIT_DRAW_BOLT = 8'd118,
				 COND_DRAW_BOLT = 8'd119,
				 DRAW_BOLT = 8'd120,
				 BITCOND_DRAW_BOLT = 8'd121,
				 INCX_DRAW_BOLT = 8'd122,
				 INCY_DRAW_BOLT = 8'd123,
				 DEC_COUNTER_DRAW_BOLT = 8'd124,
				 EXIT_DRAW_BOLT = 8'd125,
				 
				 START_DRAW_BOMB = 8'd126,
				 INIT_DRAW_BOMB = 8'd127,
				 COND_DRAW_BOMB = 8'd128,
				 DRAW_BOMB = 8'd129,
				 BITCOND_DRAW_BOMB = 8'd130,
				 INCX_DRAW_BOMB = 8'd131,
				 INCY_DRAW_BOMB = 8'd132,
				 DEC_COUNTER_DRAW_BOMB = 8'd133,
				 EXIT_DRAW_BOMB = 8'd134,
				 
				 CHECK_STATE = 8'd135,
				 
				 START_DEBOUNCE = 8'd136,
				 COND_DEBOUNCE = 8'd137,
				 INC_DEBOUNCE = 8'd138,
				 INC_LOOP = 8'd139,
				 EXIT_DEBOUNCE = 8'd140,
				 DEC_CASH = 8'd141,
				 CHECK_PRIZES = 8'd142,
				 CHECK_CASH = 8'd143,
				 
				 
				 START_DRAW_WIN = 8'd144,
				 INIT_DRAW_WIN = 8'd145,
				 COND_DRAW_WIN = 8'd146,
				 DRAW_WIN = 8'd147,
				 BITCOND_DRAW_WIN = 8'd148,
				 INCX_DRAW_WIN = 8'd149,
				 INCY_DRAW_WIN = 8'd150,
				 DEC_COUNTER_DRAW_WIN = 8'd151,
				 EXIT_DRAW_WIN = 8'd152,
				 
				 START_DRAW_LOSE = 8'd153,
				 INIT_DRAW_LOSE = 8'd154,
				 COND_DRAW_LOSE = 8'd155,
				 DRAW_LOSE = 8'd156,
				 BITCOND_DRAW_LOSE = 8'd157,
				 INCX_DRAW_LOSE = 8'd158,
				 INCY_DRAW_LOSE = 8'd159,
				 DEC_COUNTER_DRAW_LOSE = 8'd160,
				 EXIT_DRAW_LOSE = 8'd161,
				 
				 END = 8'd255;
	
	random_number rand1_mod(clk, rst, rand1);
	random_number rand2_mod(clk, rst, rand2);
	random_number rand3_mod(clk, rst, rand3);
	
	
	always @(posedge clk or negedge rst)
		if (rst == 1'b0)
			S <= START;
		else
			S <= NS;
			
	always @(*)
		case (S)
			START : 
				if (done == 1'b1)
					NS = START_DRAW_BG;
				else NS = START;
				
			START_DRAW_BG : 
			begin
				NS = INIT_DRAW_BG;
			end
			INIT_DRAW_BG : NS = COND_DRAW_BG;
			COND_DRAW_BG :
				if (backgroundImageBits[counter] == 1'b1)
					NS = DRAW_BG;
				else
					NS = BITCOND_DRAW_BG;
			
			DRAW_BG : NS = BITCOND_DRAW_BG;
			BITCOND_DRAW_BG :
				if (imageX >= backgroundImageWidth)
					NS = INCY_DRAW_BG;
				else
					NS = INCX_DRAW_BG;
					
			INCX_DRAW_BG : NS = DEC_COUNTER_DRAW_BG;
			INCY_DRAW_BG : NS = DEC_COUNTER_DRAW_BG;
			DEC_COUNTER_DRAW_BG :
				if (imageY < backgroundImageHeight)
					NS = COND_DRAW_BG;
				else
					NS = EXIT_DRAW_BG;
			
			EXIT_DRAW_BG : NS = init_left_slot;
			init_left_slot : NS = START_DRAW_START_LEFT;
			START_DRAW_START_LEFT : NS = INIT_DRAW_START_LEFT;
			INIT_DRAW_START_LEFT : NS = COND_DRAW_START_LEFT;
			COND_DRAW_START_LEFT :
				if (startImageBits[counter] == 1'b1)
					NS = DRAW_START_LEFT;
				else
					NS = BITCOND_DRAW_START_LEFT;
			
			DRAW_START_LEFT : NS = BITCOND_DRAW_START_LEFT;
			BITCOND_DRAW_START_LEFT :
				if (imageX >= startImageWidth)
					NS = INCY_DRAW_START_LEFT;
				else
					NS = INCX_DRAW_START_LEFT;
					
			INCX_DRAW_START_LEFT : NS = DEC_COUNTER_DRAW_START_LEFT;
			INCY_DRAW_START_LEFT : NS = DEC_COUNTER_DRAW_START_LEFT;
			DEC_COUNTER_DRAW_START_LEFT :
				if (imageY < startImageHeight)
					NS = COND_DRAW_START_LEFT;
				else
					NS = EXIT_DRAW_START_LEFT;
			
			EXIT_DRAW_START_LEFT : NS = init_mid_slot;
			init_mid_slot : NS = START_DRAW_START_MID;
			
			START_DRAW_START_MID : NS = INIT_DRAW_START_MID;
			INIT_DRAW_START_MID : NS = COND_DRAW_START_MID;
			COND_DRAW_START_MID :
				if (startImageBits[counter] == 1'b1)
					NS = DRAW_START_MID;
				else
					NS = BITCOND_DRAW_START_MID;
			
			DRAW_START_MID : NS = BITCOND_DRAW_START_MID;
			BITCOND_DRAW_START_MID :
				if (imageX >= startImageWidth)
					NS = INCY_DRAW_START_MID;
				else
					NS = INCX_DRAW_START_MID;
					
			INCX_DRAW_START_MID : NS = DEC_COUNTER_DRAW_START_MID;
			INCY_DRAW_START_MID : NS = DEC_COUNTER_DRAW_START_MID;
			DEC_COUNTER_DRAW_START_MID :
				if (imageY < startImageHeight)
					NS = COND_DRAW_START_MID;
				else
					NS = EXIT_DRAW_START_MID;
			
			EXIT_DRAW_START_MID : NS = init_right_slot;
			init_right_slot : NS = START_DRAW_START_RIGHT;
			START_DRAW_START_RIGHT : NS = INIT_DRAW_START_RIGHT;
			INIT_DRAW_START_RIGHT : NS = COND_DRAW_START_RIGHT;
			COND_DRAW_START_RIGHT :
				if (startImageBits[counter] == 1'b1)
					NS = DRAW_START_RIGHT;
				else
					NS = BITCOND_DRAW_START_RIGHT;
			
			DRAW_START_RIGHT : NS = BITCOND_DRAW_START_RIGHT;
			BITCOND_DRAW_START_RIGHT :
				if (imageX >= startImageWidth)
					NS = INCY_DRAW_START_RIGHT;
				else
					NS = INCX_DRAW_START_RIGHT;
					
			INCX_DRAW_START_RIGHT : NS = DEC_COUNTER_DRAW_START_RIGHT;
			INCY_DRAW_START_RIGHT : NS = DEC_COUNTER_DRAW_START_RIGHT;
			DEC_COUNTER_DRAW_START_RIGHT :
				if (imageY < startImageHeight)
					NS = COND_DRAW_START_RIGHT;
				else
					NS = EXIT_DRAW_START_RIGHT;
			
			EXIT_DRAW_START_RIGHT : NS = WAIT_FOR_INPUT;
			
			WAIT_FOR_INPUT :
				if (button[0] == 1'b0 && spinReady == 1'b1)
					NS = CLEAR_SLOTS;
				else
					NS = WAIT_FOR_INPUT;
					
			CLEAR_SLOTS : NS = START_CLEAR_LEFT;
			START_CLEAR_LEFT : NS = INIT_CLEAR_LEFT;
			INIT_CLEAR_LEFT : NS = COND_CLEAR_LEFT;
			COND_CLEAR_LEFT :
				if (clearImageBits[counter] == 1'b1)
					NS = CLEAR_LEFT;
				else
					NS = BITCOND_CLEAR_LEFT;
			
			CLEAR_LEFT : NS = BITCOND_CLEAR_LEFT;
			BITCOND_CLEAR_LEFT :
				if (imageX >= clearImageWidth)
					NS = INCY_CLEAR_LEFT;
				else
					NS = INCX_CLEAR_LEFT;
					
			INCX_CLEAR_LEFT : NS = DEC_COUNTER_CLEAR_LEFT;
			INCY_CLEAR_LEFT : NS = DEC_COUNTER_CLEAR_LEFT;
			DEC_COUNTER_CLEAR_LEFT :
				if (imageY < clearImageHeight)
					NS = COND_CLEAR_LEFT;
				else
					NS = EXIT_CLEAR_LEFT;
			
			EXIT_CLEAR_LEFT : NS = START_CLEAR_MID;
			
			
			START_CLEAR_MID : NS = INIT_CLEAR_MID;
			INIT_CLEAR_MID : NS = COND_CLEAR_MID;
			COND_CLEAR_MID :
				if (clearImageBits[counter] == 1'b1)
					NS = CLEAR_MID;
				else
					NS = BITCOND_CLEAR_MID;
			
			CLEAR_MID : NS = BITCOND_CLEAR_MID;
			BITCOND_CLEAR_MID :
				if (imageX >= clearImageWidth)
					NS = INCY_CLEAR_MID;
				else
					NS = INCX_CLEAR_MID;
					
			INCX_CLEAR_MID : NS = DEC_COUNTER_CLEAR_MID;
			INCY_CLEAR_MID : NS = DEC_COUNTER_CLEAR_MID;
			DEC_COUNTER_CLEAR_MID :
				if (imageY < clearImageHeight)
					NS = COND_CLEAR_MID;
				else
					NS = EXIT_CLEAR_MID;
			
			EXIT_CLEAR_MID : NS = START_CLEAR_RIGHT;
			
			
			START_CLEAR_RIGHT : NS = INIT_CLEAR_RIGHT;
			INIT_CLEAR_RIGHT : NS = COND_CLEAR_RIGHT;
			COND_CLEAR_RIGHT :
				if (clearImageBits[counter] == 1'b1)
					NS = CLEAR_RIGHT;
				else
					NS = BITCOND_CLEAR_RIGHT;
			
			CLEAR_RIGHT : NS = BITCOND_CLEAR_RIGHT;
			BITCOND_CLEAR_RIGHT :
				if (imageX >= clearImageWidth)
					NS = INCY_CLEAR_RIGHT;
				else
					NS = INCX_CLEAR_RIGHT;
					
			INCX_CLEAR_RIGHT : NS = DEC_COUNTER_CLEAR_RIGHT;
			INCY_CLEAR_RIGHT : NS = DEC_COUNTER_CLEAR_RIGHT;
			DEC_COUNTER_CLEAR_RIGHT :
				if (imageY < clearImageHeight)
					NS = COND_CLEAR_RIGHT;
				else
					NS = EXIT_CLEAR_RIGHT;
			
			EXIT_CLEAR_RIGHT : NS = CHECK_SLOT1;
			CHECK_SLOT1 :
				case (rand1)
					3'd0 : NS = START_DRAW_SEVEN;
					3'd1 : NS = START_DRAW_ORANGE;
					3'd2 : NS = START_DRAW_LEMON;
					3'd3 : NS = START_DRAW_COIN;
					3'd4 : NS = START_DRAW_DOLLAR;
					3'd5 : NS = START_DRAW_BOLT;
					default : NS = START_DRAW_BOMB;
				endcase
			
			CHECK_SLOT2 :
				case (rand2)
					3'd0 : NS = START_DRAW_SEVEN;
					3'd1 : NS = START_DRAW_ORANGE;
					3'd2 : NS = START_DRAW_LEMON;
					3'd3 : NS = START_DRAW_COIN;
					3'd4 : NS = START_DRAW_DOLLAR;
					3'd5 : NS = START_DRAW_BOLT;
					default : NS = START_DRAW_BOMB;
				endcase
			
			CHECK_SLOT3 :
				case (rand3)
					3'd0 : NS = START_DRAW_SEVEN;
					3'd1 : NS = START_DRAW_ORANGE;
					3'd2 : NS = START_DRAW_LEMON;
					3'd3 : NS = START_DRAW_COIN;
					3'd4 : NS = START_DRAW_DOLLAR;
					3'd5 : NS = START_DRAW_BOLT;
					default : NS = START_DRAW_BOMB;
				endcase

			CHECK_STATE :
				case (currentCheckState)
					2'd0 : NS = CHECK_SLOT1;
					2'd1 : NS = CHECK_SLOT2;
					2'd2 : NS = CHECK_SLOT3;
					2'd3 : NS = START_DEBOUNCE;
					default : begin end
				endcase
				
			START_DEBOUNCE : NS = COND_DEBOUNCE;
			COND_DEBOUNCE : 
				if (loopCounter >= 4'd7)
					NS = EXIT_DEBOUNCE;
				else if (debounceCounter >= 26'd5000000)
					NS = INC_LOOP;
				else
					NS = INC_DEBOUNCE;
					
			INC_LOOP : NS = CLEAR_SLOTS;
			
			INC_DEBOUNCE : NS = COND_DEBOUNCE;
			EXIT_DEBOUNCE : NS = DEC_CASH;
			DEC_CASH : NS = CHECK_PRIZES;
			
			CHECK_PRIZES : NS = CHECK_CASH;

			CHECK_CASH :
				if (player_balance >= 7'd100)
					NS = START_DRAW_WIN;
				else if (player_balance < 3'd5)
					NS = START_DRAW_LOSE;
				else
					NS = WAIT_FOR_INPUT;
			
			
			START_DRAW_WIN : NS = INIT_DRAW_WIN;
			INIT_DRAW_WIN : NS = COND_DRAW_WIN;
			COND_DRAW_WIN :
				if (winImageBits[counter] == 1'b1)
					NS = DRAW_WIN;
				else
					NS = BITCOND_DRAW_WIN;
			
			DRAW_WIN : NS = BITCOND_DRAW_WIN;
			BITCOND_DRAW_WIN :
				if (imageX >= winImageWidth)
					NS = INCY_DRAW_WIN;
				else
					NS = INCX_DRAW_WIN;
					
			INCX_DRAW_WIN : NS = DEC_COUNTER_DRAW_WIN;
			INCY_DRAW_WIN : NS = DEC_COUNTER_DRAW_WIN;
			DEC_COUNTER_DRAW_WIN :
				if (imageY < winImageHeight)
					NS = COND_DRAW_WIN;
				else
					NS = EXIT_DRAW_WIN;
			
			EXIT_DRAW_WIN : NS = END;
			
			
			START_DRAW_LOSE : NS = INIT_DRAW_LOSE;
			INIT_DRAW_LOSE : NS = COND_DRAW_LOSE;
			COND_DRAW_LOSE :
				if (loseImageBits[counter] == 1'b1)
					NS = DRAW_LOSE;
				else
					NS = BITCOND_DRAW_LOSE;
			
			DRAW_LOSE : NS = BITCOND_DRAW_LOSE;
			BITCOND_DRAW_LOSE :
				if (imageX >= loseImageWidth)
					NS = INCY_DRAW_LOSE;
				else
					NS = INCX_DRAW_LOSE;
					
			INCX_DRAW_LOSE : NS = DEC_COUNTER_DRAW_LOSE;
			INCY_DRAW_LOSE : NS = DEC_COUNTER_DRAW_LOSE;
			DEC_COUNTER_DRAW_LOSE :
				if (imageY < loseImageHeight)
					NS = COND_DRAW_LOSE;
				else
					NS = EXIT_DRAW_LOSE;
			
			EXIT_DRAW_LOSE : NS = END;
			
				
			START_DRAW_SEVEN : NS = INIT_DRAW_SEVEN;
			INIT_DRAW_SEVEN : NS = COND_DRAW_SEVEN;
			COND_DRAW_SEVEN :
				if (sevenImageBits[counter] == 1'b1)
					NS = DRAW_SEVEN;
				else
					NS = BITCOND_DRAW_SEVEN;
			
			DRAW_SEVEN : NS = BITCOND_DRAW_SEVEN;
			BITCOND_DRAW_SEVEN :
				if (imageX >= sevenImageWidth)
					NS = INCY_DRAW_SEVEN;
				else
					NS = INCX_DRAW_SEVEN;
					
			INCX_DRAW_SEVEN : NS = DEC_COUNTER_DRAW_SEVEN;
			INCY_DRAW_SEVEN : NS = DEC_COUNTER_DRAW_SEVEN;
			DEC_COUNTER_DRAW_SEVEN :
				if (imageY < sevenImageHeight)
					NS = COND_DRAW_SEVEN;
				else
					NS = EXIT_DRAW_SEVEN;
			
			EXIT_DRAW_SEVEN : NS = CHECK_STATE;
			
			START_DRAW_ORANGE : NS = INIT_DRAW_ORANGE;
			INIT_DRAW_ORANGE : NS = COND_DRAW_ORANGE;
			COND_DRAW_ORANGE :
				if (orangeImageBits[counter] == 1'b1)
					NS = DRAW_ORANGE;
				else
					NS = BITCOND_DRAW_ORANGE;
			
			DRAW_ORANGE : NS = BITCOND_DRAW_ORANGE;
			BITCOND_DRAW_ORANGE :
				if (imageX >= orangeImageWidth)
					NS = INCY_DRAW_ORANGE;
				else
					NS = INCX_DRAW_ORANGE;
					
			INCX_DRAW_ORANGE : NS = DEC_COUNTER_DRAW_ORANGE;
			INCY_DRAW_ORANGE : NS = DEC_COUNTER_DRAW_ORANGE;
			DEC_COUNTER_DRAW_ORANGE :
				if (imageY < orangeImageHeight)
					NS = COND_DRAW_ORANGE;
				else
					NS = EXIT_DRAW_ORANGE;
			
			EXIT_DRAW_ORANGE : NS = CHECK_STATE;
			
			
			START_DRAW_LEMON : NS = INIT_DRAW_LEMON;
			INIT_DRAW_LEMON : NS = COND_DRAW_LEMON;
			COND_DRAW_LEMON :
				if (lemonImageBits[counter] == 1'b1)
					NS = DRAW_LEMON;
				else
					NS = BITCOND_DRAW_LEMON;
			
			DRAW_LEMON : NS = BITCOND_DRAW_LEMON;
			BITCOND_DRAW_LEMON :
				if (imageX >= lemonImageWidth)
					NS = INCY_DRAW_LEMON;
				else
					NS = INCX_DRAW_LEMON;
					
			INCX_DRAW_LEMON : NS = DEC_COUNTER_DRAW_LEMON;
			INCY_DRAW_LEMON : NS = DEC_COUNTER_DRAW_LEMON;
			DEC_COUNTER_DRAW_LEMON :
				if (imageY < lemonImageHeight)
					NS = COND_DRAW_LEMON;
				else
					NS = EXIT_DRAW_LEMON;
			
			EXIT_DRAW_LEMON : NS = CHECK_STATE;
			
			
			START_DRAW_COIN : NS = INIT_DRAW_COIN;
			INIT_DRAW_COIN : NS = COND_DRAW_COIN;
			COND_DRAW_COIN :
				if (coinImageBits[counter] == 1'b1)
					NS = DRAW_COIN;
				else
					NS = BITCOND_DRAW_COIN;
			
			DRAW_COIN : NS = BITCOND_DRAW_COIN;
			BITCOND_DRAW_COIN :
				if (imageX >= coinImageWidth)
					NS = INCY_DRAW_COIN;
				else
					NS = INCX_DRAW_COIN;
					
			INCX_DRAW_COIN : NS = DEC_COUNTER_DRAW_COIN;
			INCY_DRAW_COIN : NS = DEC_COUNTER_DRAW_COIN;
			DEC_COUNTER_DRAW_COIN :
				if (imageY < coinImageHeight)
					NS = COND_DRAW_COIN;
				else
					NS = EXIT_DRAW_COIN;
			
			EXIT_DRAW_COIN : NS = CHECK_STATE;
			
			
			START_DRAW_DOLLAR : NS = INIT_DRAW_DOLLAR;
			INIT_DRAW_DOLLAR : NS = COND_DRAW_DOLLAR;
			COND_DRAW_DOLLAR :
				if (dollarImageBits[counter] == 1'b1)
					NS = DRAW_DOLLAR;
				else
					NS = BITCOND_DRAW_DOLLAR;
			
			DRAW_DOLLAR : NS = BITCOND_DRAW_DOLLAR;
			BITCOND_DRAW_DOLLAR :
				if (imageX >= dollarImageWidth)
					NS = INCY_DRAW_DOLLAR;
				else
					NS = INCX_DRAW_DOLLAR;
					
			INCX_DRAW_DOLLAR : NS = DEC_COUNTER_DRAW_DOLLAR;
			INCY_DRAW_DOLLAR : NS = DEC_COUNTER_DRAW_DOLLAR;
			DEC_COUNTER_DRAW_DOLLAR :
				if (imageY < dollarImageHeight)
					NS = COND_DRAW_DOLLAR;
				else
					NS = EXIT_DRAW_DOLLAR;
			
			EXIT_DRAW_DOLLAR : NS = CHECK_STATE;
			
			
			START_DRAW_BOLT : NS = INIT_DRAW_BOLT;
			INIT_DRAW_BOLT : NS = COND_DRAW_BOLT;
			COND_DRAW_BOLT :
				if (boltImageBits[counter] == 1'b1)
					NS = DRAW_BOLT;
				else
					NS = BITCOND_DRAW_BOLT;
			
			DRAW_BOLT : NS = BITCOND_DRAW_BOLT;
			BITCOND_DRAW_BOLT :
				if (imageX >= boltImageWidth)
					NS = INCY_DRAW_BOLT;
				else
					NS = INCX_DRAW_BOLT;
					
			INCX_DRAW_BOLT : NS = DEC_COUNTER_DRAW_BOLT;
			INCY_DRAW_BOLT : NS = DEC_COUNTER_DRAW_BOLT;
			DEC_COUNTER_DRAW_BOLT :
				if (imageY < boltImageHeight)
					NS = COND_DRAW_BOLT;
				else
					NS = EXIT_DRAW_BOLT;
			
			EXIT_DRAW_BOLT : NS = CHECK_STATE;
			
			
			START_DRAW_BOMB : NS = INIT_DRAW_BOMB;
			INIT_DRAW_BOMB : NS = COND_DRAW_BOMB;
			COND_DRAW_BOMB :
				if (bombImageBits[counter] == 1'b1)
					NS = DRAW_BOMB;
				else
					NS = BITCOND_DRAW_BOMB;
			
			DRAW_BOMB : NS = BITCOND_DRAW_BOMB;
			BITCOND_DRAW_BOMB :
				if (imageX >= bombImageWidth)
					NS = INCY_DRAW_BOMB;
				else
					NS = INCX_DRAW_BOMB;
					
			INCX_DRAW_BOMB : NS = DEC_COUNTER_DRAW_BOMB;
			INCY_DRAW_BOMB : NS = DEC_COUNTER_DRAW_BOMB;
			DEC_COUNTER_DRAW_BOMB :
				if (imageY < bombImageHeight)
					NS = COND_DRAW_BOMB;
				else
					NS = EXIT_DRAW_BOMB;
			
			EXIT_DRAW_BOMB : NS = CHECK_STATE;
			
				
			END : NS = END;
			
		endcase
			
			
	always @(posedge clk or negedge rst)
		if (rst == 1'b0)
		begin
			currentInitX <= 64'b0;
			done <= 1'b0;
			colour <= 6'b000000;
			x <= 8'b00000000;
			y <= 8'b00000000;
			draw <= 18'b0;
			light1 <= 1'b0;
			light2 <= 1'b0;
			imageX <= 64'b0;
			imageY <= 64'b0;
			counter <= 64'b0;
			currentCheckState <= 2'd0;
			spinReady <= 1'b1;
			debounceCounter <= 64'b0;
			player_balance <= 10'd50;
			currentLeftSlot <= 3'd0;
			currentMidSlot <= 3'd0;
			currentRightSlot <= 3'd0;
		end
		else
			case (S)
				START :
					if (draw < 17'b10000000000000000)
					begin
						done <= 1'b0;
						x <= draw[7:0];
						y <= draw[16:8];
						draw <= draw + 1'b1;
						colour <= 6'b111111;
					end
					else
					begin
						done <= 1'b1;
						draw <= 17'b0;
					end

				START_DRAW_BG : begin end
				INIT_DRAW_BG : counter <= backgroundImageStart;
				COND_DRAW_BG : begin end
				DRAW_BG :
				begin
					colour <= 6'b110000;
					x <= initXBG + imageX;
					y <= initYBG + imageY;
				end
				
				BITCOND_DRAW_BG : begin end
				INCX_DRAW_BG : imageX <= imageX + 1'b1;
				INCY_DRAW_BG :
				begin
					imageX <= 64'b0;
					imageY <= imageY + 1'b1;
				end
				DEC_COUNTER_DRAW_BG : counter <= counter - 1'b1;
				EXIT_DRAW_BG :
				begin
					imageX <= 64'b0;
					imageY <= 64'b0;
				end
					
				init_left_slot : begin end
				START_DRAW_START_LEFT : begin end
				INIT_DRAW_START_LEFT : counter <= startImageStart;
				COND_DRAW_START_LEFT : begin end
				DRAW_START_LEFT :
				begin
					colour <= 6'b001100;
					x <= initXStartLeftSlot + imageX;
					y <= initYStartLeftSlot + imageY;
				end
				
				BITCOND_DRAW_START_LEFT : begin end
				INCX_DRAW_START_LEFT : imageX <= imageX + 1'b1;
				INCY_DRAW_START_LEFT :
				begin
					imageX <= 64'b0;
					imageY <= imageY + 1'b1;
				end
				DEC_COUNTER_DRAW_START_LEFT : counter <= counter - 1'b1;
				EXIT_DRAW_START_LEFT :
				begin
					imageX <= 64'b0;
					imageY <= 64'b0;
				end
				
				init_mid_slot : begin end
				START_DRAW_START_MID : begin end
				INIT_DRAW_START_MID : counter <= startImageStart;
				COND_DRAW_START_MID : begin end
				DRAW_START_MID :
				begin
					colour <= 6'b001100;
					x <= initXStartMidSlot + imageX;
					y <= initYStartMidSlot + imageY;
				end
				
				BITCOND_DRAW_START_MID : begin end
				INCX_DRAW_START_MID : imageX <= imageX + 1'b1;
				INCY_DRAW_START_MID :
				begin
					imageX <= 64'b0;
					imageY <= imageY + 1'b1;
				end
				DEC_COUNTER_DRAW_START_MID : counter <= counter - 1'b1;
				EXIT_DRAW_START_MID :
				begin
					imageX <= 64'b0;
					imageY <= 64'b0;
				end
				
				init_right_slot : begin end
				START_DRAW_START_RIGHT : begin end
				INIT_DRAW_START_RIGHT : counter <= startImageStart;
				COND_DRAW_START_RIGHT : begin end
				DRAW_START_RIGHT :
				begin
					colour <= 6'b001100;
					x <= initXStartRightSlot + imageX;
					y <= initYStartRightSlot + imageY;
				end
				
				BITCOND_DRAW_START_RIGHT : begin end
				INCX_DRAW_START_RIGHT : imageX <= imageX + 1'b1;
				INCY_DRAW_START_RIGHT :
				begin
					imageX <= 64'b0;
					imageY <= imageY + 1'b1;
				end
				DEC_COUNTER_DRAW_START_RIGHT : counter <= counter - 1'b1;
				EXIT_DRAW_START_RIGHT :
				begin
					imageX <= 64'b0;
					imageY <= 64'b0;
				end
				
				START_DEBOUNCE : begin debounceCounter <= 64'b0; end
				COND_DEBOUNCE : begin end
				INC_DEBOUNCE : debounceCounter <= debounceCounter + 1'b1;
				INC_LOOP :
				begin
					debounceCounter <= 64'b0;
					loopCounter <= loopCounter + 1'b1;
				end
				EXIT_DEBOUNCE :
				begin
					loopCounter <= 4'd0;
					spinReady <= 1'b1;
				end
				
				DEC_CASH : player_balance <= player_balance - 3'd5;
				
				CHECK_PRIZES :
				begin
					if (currentLeftSlot == currentMidSlot && currentMidSlot == currentRightSlot)
						case (currentMidSlot)
							3'd0 : player_balance <= player_balance + 4'd5;
							3'd1 : player_balance <= player_balance + 5'd10;
							3'd2 : player_balance <= player_balance + 6'd25;
							3'd3 : player_balance <= player_balance + 7'd50;
							3'd4 : player_balance <= player_balance + 7'd75;
							3'd5 : player_balance <= 7'd100;
							default : player_balance <= 10'd0;
						endcase
				end
				
				WAIT_FOR_INPUT :
				begin
					light2 <= 1'b1;
					currentCheckState <= 2'd0;
				end

				CLEAR_SLOTS : begin spinReady <= 1'b0; light2 <= 1'b0; end

				START_CLEAR_LEFT : begin end
				INIT_CLEAR_LEFT : counter <= clearImageStart;
				COND_CLEAR_LEFT : begin end
				CLEAR_LEFT :
				begin
					colour <= 6'b111111;
					x <= initXStartLeftSlot + imageX;
					y <= initYStartLeftSlot + imageY;
				end
				
				BITCOND_CLEAR_LEFT : begin end
				INCX_CLEAR_LEFT : imageX <= imageX + 1'b1;
				INCY_CLEAR_LEFT :
				begin
					imageX <= 64'b0;
					imageY <= imageY + 1'b1;
				end
				DEC_COUNTER_CLEAR_LEFT : counter <= counter - 1'b1;
				EXIT_CLEAR_LEFT :
				begin
					imageX <= 64'b0;
					imageY <= 64'b0;
				end
				
				START_CLEAR_MID : begin end
				INIT_CLEAR_MID : counter <= clearImageStart;
				COND_CLEAR_MID : begin end
				CLEAR_MID :
				begin
					colour <= 6'b111111;
					x <= initXStartMidSlot + imageX;
					y <= initYStartMidSlot + imageY;
				end
				
				BITCOND_CLEAR_MID : begin end
				INCX_CLEAR_MID : imageX <= imageX + 1'b1;
				INCY_CLEAR_MID :
				begin
					imageX <= 64'b0;
					imageY <= imageY + 1'b1;
				end
				DEC_COUNTER_CLEAR_MID : counter <= counter - 1'b1;
				EXIT_CLEAR_MID :
				begin
					imageX <= 64'b0;
					imageY <= 64'b0;
				end
				
				START_CLEAR_RIGHT : begin end
				INIT_CLEAR_RIGHT : counter <= clearImageStart;
				COND_CLEAR_RIGHT : begin end
				CLEAR_RIGHT :
				begin
					colour <= 6'b111111;
					x <= initXStartRightSlot + imageX;
					y <= initYStartRightSlot + imageY;
				end
				
				BITCOND_CLEAR_RIGHT : begin end
				INCX_CLEAR_RIGHT : imageX <= imageX + 1'b1;
				INCY_CLEAR_RIGHT :
				begin
					imageX <= 64'b0;
					imageY <= imageY + 1'b1;
				end
				DEC_COUNTER_CLEAR_RIGHT : counter <= counter - 1'b1;
				EXIT_CLEAR_RIGHT :
				begin
					imageX <= 64'b0;
					imageY <= 64'b0;
				end
				
				CHECK_SLOT1 :
				begin
					currentCheckState <= 2'd1;
					currentInitX <= initXStartLeftSlot;
				end
				CHECK_SLOT2 :
				begin
					currentCheckState <= 2'd2;
					currentInitX <= initXStartMidSlot;
				end
				CHECK_SLOT3 :
				begin
					currentCheckState <= 2'd3;
					currentInitX <= initXStartRightSlot;
				end
				
				START_DRAW_SEVEN : begin end
				INIT_DRAW_SEVEN : counter <= sevenImageStart;
				COND_DRAW_SEVEN : begin end
				DRAW_SEVEN :
				begin
					colour <= 6'b110000;
					x <= currentInitX + imageX;
					y <= initYStartLeftSlot + imageY;
				end
				
				BITCOND_DRAW_SEVEN : begin end
				INCX_DRAW_SEVEN : imageX <= imageX + 1'b1;
				INCY_DRAW_SEVEN :
				begin
					imageX <= 64'b0;
					imageY <= imageY + 1'b1;
				end
				DEC_COUNTER_DRAW_SEVEN : counter <= counter - 1'b1;
				EXIT_DRAW_SEVEN :
				begin
					imageX <= 64'b0;
					imageY <= 64'b0;
					case (currentInitX)
						initXStartLeftSlot : currentLeftSlot <= 3'd0;
						initXStartMidSlot : currentMidSlot <= 3'd0;
						initXStartRightSlot : currentRightSlot <= 3'd0;
						default : begin end
					endcase
				end
				
				START_DRAW_ORANGE : begin end
				INIT_DRAW_ORANGE : counter <= orangeImageStart;
				COND_DRAW_ORANGE : begin end
				DRAW_ORANGE :
				begin
					colour <= 6'b111000;
					x <= currentInitX + imageX;
					y <= initYStartLeftSlot + imageY;
				end
				
				BITCOND_DRAW_ORANGE : begin end
				INCX_DRAW_ORANGE : imageX <= imageX + 1'b1;
				INCY_DRAW_ORANGE :
				begin
					imageX <= 64'b0;
					imageY <= imageY + 1'b1;
				end
				DEC_COUNTER_DRAW_ORANGE : counter <= counter - 1'b1;
				EXIT_DRAW_ORANGE :
				begin
					imageX <= 64'b0;
					imageY <= 64'b0;
					case (currentInitX)
						initXStartLeftSlot : currentLeftSlot <= 3'd1;
						initXStartMidSlot : currentMidSlot <= 3'd1;
						initXStartRightSlot : currentRightSlot <= 3'd1;
						default : begin end
					endcase
				end
				
				START_DRAW_LEMON : begin end
				INIT_DRAW_LEMON : counter <= lemonImageStart;
				COND_DRAW_LEMON : begin end
				DRAW_LEMON :
				begin
					colour <= 6'b111100;
					x <= currentInitX + imageX;
					y <= initYStartLeftSlot + imageY;
				end
				
				BITCOND_DRAW_LEMON : begin end
				INCX_DRAW_LEMON : imageX <= imageX + 1'b1;
				INCY_DRAW_LEMON :
				begin
					imageX <= 64'b0;
					imageY <= imageY + 1'b1;
				end
				DEC_COUNTER_DRAW_LEMON : counter <= counter - 1'b1;
				EXIT_DRAW_LEMON :
				begin
					imageX <= 64'b0;
					imageY <= 64'b0;
					case (currentInitX)
						initXStartLeftSlot : currentLeftSlot <= 3'd2;
						initXStartMidSlot : currentMidSlot <= 3'd2;
						initXStartRightSlot : currentRightSlot <= 3'd2;
						default : begin end
					endcase
				end
				
				START_DRAW_COIN : begin end
				INIT_DRAW_COIN : counter <= coinImageStart;
				COND_DRAW_COIN : begin end
				DRAW_COIN :
				begin
					colour <= 6'b101000;
					x <= currentInitX + imageX;
					y <= initYStartLeftSlot + imageY;
				end
				
				BITCOND_DRAW_COIN : begin end
				INCX_DRAW_COIN : imageX <= imageX + 1'b1;
				INCY_DRAW_COIN :
				begin
					imageX <= 64'b0;
					imageY <= imageY + 1'b1;
				end
				DEC_COUNTER_DRAW_COIN : counter <= counter - 1'b1;
				EXIT_DRAW_COIN :
				begin
					imageX <= 64'b0;
					imageY <= 64'b0;
					case (currentInitX)
						initXStartLeftSlot : currentLeftSlot <= 3'd3;
						initXStartMidSlot : currentMidSlot <= 3'd3;
						initXStartRightSlot : currentRightSlot <= 3'd3;
						default : begin end
					endcase
				end
				
				START_DRAW_DOLLAR : begin end
				INIT_DRAW_DOLLAR : counter <= dollarImageStart;
				COND_DRAW_DOLLAR : begin end
				DRAW_DOLLAR :
				begin
					colour <= 6'b001100;
					x <= currentInitX + imageX;
					y <= initYStartLeftSlot + imageY;
				end
				
				BITCOND_DRAW_DOLLAR : begin end
				INCX_DRAW_DOLLAR : imageX <= imageX + 1'b1;
				INCY_DRAW_DOLLAR :
				begin
					imageX <= 64'b0;
					imageY <= imageY + 1'b1;
				end
				DEC_COUNTER_DRAW_DOLLAR : counter <= counter - 1'b1;
				EXIT_DRAW_DOLLAR :
				begin
					imageX <= 64'b0;
					imageY <= 64'b0;
					case (currentInitX)
						initXStartLeftSlot : currentLeftSlot <= 3'd4;
						initXStartMidSlot : currentMidSlot <= 3'd4;
						initXStartRightSlot : currentRightSlot <= 3'd4;
						default : begin end
					endcase
				end
				
				START_DRAW_BOLT : begin end
				INIT_DRAW_BOLT : counter <= boltImageStart;
				COND_DRAW_BOLT : begin end
				DRAW_BOLT :
				begin
					colour <= 6'b111100;
					x <= currentInitX + imageX;
					y <= initYStartLeftSlot + imageY;
				end
				
				BITCOND_DRAW_BOLT : begin end
				INCX_DRAW_BOLT : imageX <= imageX + 1'b1;
				INCY_DRAW_BOLT :
				begin
					imageX <= 64'b0;
					imageY <= imageY + 1'b1;
				end
				DEC_COUNTER_DRAW_BOLT : counter <= counter - 1'b1;
				EXIT_DRAW_BOLT :
				begin
					imageX <= 64'b0;
					imageY <= 64'b0;
					case (currentInitX)
						initXStartLeftSlot : currentLeftSlot <= 3'd5;
						initXStartMidSlot : currentMidSlot <= 3'd5;
						initXStartRightSlot : currentRightSlot <= 3'd5;
						default : begin end
					endcase
				end
				
				START_DRAW_BOMB : begin end
				INIT_DRAW_BOMB : counter <= bombImageStart;
				COND_DRAW_BOMB : begin end
				DRAW_BOMB :
				begin
					colour <= 6'b000000;
					x <= currentInitX + imageX;
					y <= initYStartLeftSlot + imageY;
				end
				
				BITCOND_DRAW_BOMB : begin end
				INCX_DRAW_BOMB : imageX <= imageX + 1'b1;
				INCY_DRAW_BOMB :
				begin
					imageX <= 64'b0;
					imageY <= imageY + 1'b1;
				end
				DEC_COUNTER_DRAW_BOMB : counter <= counter - 1'b1;
				EXIT_DRAW_BOMB :
				begin
					imageX <= 64'b0;
					imageY <= 64'b0;
					case (currentInitX)
						initXStartLeftSlot : currentLeftSlot <= 3'd6;
						initXStartMidSlot : currentMidSlot <= 3'd6;
						initXStartRightSlot : currentRightSlot <= 3'd6;
						default : begin end
					endcase
				end
				
				START_DRAW_WIN : begin end
				INIT_DRAW_WIN : counter <= winImageStart;
				COND_DRAW_WIN : begin end
				DRAW_WIN :
				begin
					colour <= 6'b110000;
					x <= initXEnd + imageX;
					y <= initYEnd + imageY;
				end
				
				BITCOND_DRAW_WIN : begin end
				INCX_DRAW_WIN : imageX <= imageX + 1'b1;
				INCY_DRAW_WIN :
				begin
					imageX <= 64'b0;
					imageY <= imageY + 1'b1;
				end
				DEC_COUNTER_DRAW_WIN : counter <= counter - 1'b1;
				EXIT_DRAW_WIN :
				begin
					imageX <= 64'b0;
					imageY <= 64'b0;
				end
				
				END : done <= 1'b1;
				
				
				START_DRAW_LOSE : begin end
				INIT_DRAW_LOSE : counter <= loseImageStart;
				COND_DRAW_LOSE : begin end
				DRAW_LOSE :
				begin
					colour <= 6'b110000;
					x <= initXEnd + imageX;
					y <= initYEnd + imageY;
				end
				
				BITCOND_DRAW_LOSE : begin end
				INCX_DRAW_LOSE : imageX <= imageX + 1'b1;
				INCY_DRAW_LOSE :
				begin
					imageX <= 64'b0;
					imageY <= imageY + 1'b1;
				end
				DEC_COUNTER_DRAW_LOSE : counter <= counter - 1'b1;
				EXIT_DRAW_LOSE :
				begin
					imageX <= 64'b0;
					imageY <= 64'b0;
				end
				
				END : done <= 1'b1;
			endcase
	
endmodule 


module clock (input clock, output clk);
	reg [19:0] frame_counter;
	reg frame;

	always@(posedge clock)
	  begin
		 if (frame_counter == 20'b0) begin
			frame_counter = 20'd833332;  // This divisor gives us ~60 frames per second
			frame = 1'b1;
		 end 
		 
		 else 
		 begin
			frame_counter = frame_counter - 1'b1;
			frame = 1'b0;
		 end
	  end

	assign clk = frame;
endmodule
